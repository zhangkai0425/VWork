module int_mnt();

endmodule
