
`timescale 1ns/100ps

`define CLK_PERIOD          10
`define TCLK_PERIOD         40
`define MAX_RUN_TIME        32'h3000000

`define SOC_TOP             tb.x_soc
//`define RTL_MEM             tb.x_soc.x_aqe_iram.x_f_spsram_large
`define CPU_TOP             tb.x_soc.x_cpu_sub_system
`define tb_retire0          `CPU_TOP.core0_pad_retire0
`define retire0_pc          `CPU_TOP.core0_pad_retire0_pc[39:0]
`define tb_retire1          `CPU_TOP.core0_pad_retire1
`define retire1_pc          `CPU_TOP.core0_pad_retire1_pc[39:0]
`define CPU_CLK             `CPU_TOP.pll_cpu_clk
`define CPU_RST             `CPU_TOP.pad_cpu_rst_b
`define clk_en              `CPU_TOP.axim_clk_en

// `define APB_BASE_ADDR       40'h4000000000
`define APB_BASE_ADDR       40'hb0000000

module tb();
  reg clk;
  reg rst_b;

  integer FILE;
  
  initial
  begin
    clk =0;
    forever begin
      #(`CLK_PERIOD/2) clk = ~clk;
    end
  end
  
  initial
  begin
    rst_b = 1;
    #100;
    rst_b = 0;
    #100;
    rst_b = 1;
  end
  
  // test dual port:
  reg uart2sys_en;
  reg [39:0] uart2sys_addr;
  reg [127:0] uart2sys_data;
  reg sys_wren;
  reg [39:0] sys_final_addr;
  reg [127:0] sys_data;
  initial
  begin
    uart2sys_en = 0;
    sys_wren = 0;
    uart2sys_addr = 40'h0002000020;
    sys_final_addr = 40'h0002000020; 
    uart2sys_data = 128'h7;
    sys_data = 128'h8;
    #(`CLK_PERIOD*2000);
    uart2sys_en = 1;
    #(`CLK_PERIOD*10);
    uart2sys_en = 0;
    #(`CLK_PERIOD*10);
    sys_wren = 1;
    #(`CLK_PERIOD*100);
    sys_wren = 0;
  end
  // test dual port end;
  integer i;
  reg [31:0] mem_inst_temp [16777216:0];
  reg [31:0] mem_data_temp [16777216:0];
  integer j;
  initial
  begin
    $display("\t********* Init Program *********");
    $display("\t********* Wipe memory to 0 *********");
//    for(i=0; i < 32'h1000000; i=i+1)
//    begin
//      `RTL_MEM.ram0.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram1.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram2.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram3.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram4.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram5.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram6.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram7.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram8.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram9.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram10.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram11.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram12.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram13.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram14.mem[i][7:0] = 8'h0;
//      `RTL_MEM.ram15.mem[i][7:0] = 8'h0;
//    end
  
    $display("\t********* Read program *********");
    $readmemh("inst.mem", mem_inst_temp);
    $readmemh("data.mem", mem_data_temp);
  
    $display("\t********* Load program to memory *********");
    i=0;
//    for(j=0;i<32'h4000;i=j/4)
//    begin
//      `RTL_MEM.ram0.mem[i][7:0] = mem_inst_temp[j][31:24];
//      `RTL_MEM.ram1.mem[i][7:0] = mem_inst_temp[j][23:16];
//      `RTL_MEM.ram2.mem[i][7:0] = mem_inst_temp[j][15: 8];
//      `RTL_MEM.ram3.mem[i][7:0] = mem_inst_temp[j][ 7: 0];
//      j = j+1;
//      `RTL_MEM.ram4.mem[i][7:0] = mem_inst_temp[j][31:24];
//      `RTL_MEM.ram5.mem[i][7:0] = mem_inst_temp[j][23:16];
//      `RTL_MEM.ram6.mem[i][7:0] = mem_inst_temp[j][15: 8];
//      `RTL_MEM.ram7.mem[i][7:0] = mem_inst_temp[j][ 7: 0];
//      j = j+1;
//      `RTL_MEM.ram8.mem[i][7:0] = mem_inst_temp[j][31:24];
//      `RTL_MEM.ram9.mem[i][7:0] = mem_inst_temp[j][23:16];
//      `RTL_MEM.ram10.mem[i][7:0] = mem_inst_temp[j][15: 8];
//      `RTL_MEM.ram11.mem[i][7:0] = mem_inst_temp[j][ 7: 0];
//      j = j+1;
//      `RTL_MEM.ram12.mem[i][7:0] = mem_inst_temp[j][31:24];
//      `RTL_MEM.ram13.mem[i][7:0] = mem_inst_temp[j][23:16];
//      `RTL_MEM.ram14.mem[i][7:0] = mem_inst_temp[j][15: 8];
//      `RTL_MEM.ram15.mem[i][7:0] = mem_inst_temp[j][ 7: 0];
//      j = j+1;
//    end
  end

  initial
  begin
  #(`MAX_RUN_TIME * `CLK_PERIOD);
    $display("**********************************************");
    $display("*   meeting max simulation time, stop!       *");
    $display("**********************************************");
    FILE = $fopen("run_case.report","w");
    $fwrite(FILE,"TEST FAIL");   
  $finish;
  end

  reg [31:0] cycle_count;
  
  `define LAST_CYCLE 50000
  always @(posedge clk or negedge rst_b)
  begin
    if(!rst_b)
      cycle_count[31:0] <= 32'b1;
    else 
      cycle_count[31:0] <= cycle_count[31:0] + 1'b1;
  end
  
  reg [31:0] cpu_awaddr;
  reg [3:0]  cpu_awlen;
  reg [15:0] cpu_wstrb;
  reg        cpu_wvalid;
  reg [63:0] value0;
  reg [63:0] value1;
  reg [63:0] value2;
  
  always @(posedge `CPU_CLK)
  begin
    cpu_awlen[3:0]   <= `SOC_TOP.x_aqe_iram.awlen[3:0];
    cpu_awaddr[31:0] <= `SOC_TOP.x_aqe_iram.mem_addr[31:0];
    cpu_wvalid       <= `SOC_TOP.biu_pad_wvalid;
    cpu_wstrb        <= `SOC_TOP.biu_pad_wstrb;
 
    value0              <= `CPU_TOP.x_C908_TOP.x_pc_top_0.x_pc_core.x_pc_iu_top.x_pc_iu_dp.dp_pipe0_ex4_wb_data[63:0];
    value1              <= `CPU_TOP.x_C908_TOP.x_pc_top_0.x_pc_core.x_pc_iu_top.x_pc_iu_dp.dp_pipe1_ex4_wb_data[63:0];
  end
  
  always @(posedge `CPU_CLK)
  begin
      if(value0 == 64'h444333222 || value1 == 64'h444333222 || value2 == 64'h444333222)
    begin
      $display("**********************************************");
      $display("*    simulation finished successfully        *");
      $display("**********************************************");
     #10;
     FILE = $fopen("run_case.report","w");
     $fwrite(FILE,"TEST PASS");   
  
     $finish;
    end
      else if (value0 == 64'h2382348720 || value1 == 64'h2382348720 || value2 == 64'h444333222)
    begin
     $display("**********************************************");
     $display("*    simulation finished with error          *");
     $display("**********************************************");
     #10;
     FILE = $fopen("run_case.report","w");
     $fwrite(FILE,"TEST FAIL");   
  
     $finish;
    end
  
    else if((cpu_awlen[3:0] == 4'b0) &&
       (cpu_awaddr[31:0] == 32'h01ff_fff0) &&
        cpu_wvalid &&
       `clk_en)
    begin
     if(cpu_wstrb[15:0] == 16'hf)
     begin
        $write("%c", `SOC_TOP.biu_pad_wdata[7:0]);
     end
     else if(cpu_wstrb[15:0] == 16'hf0)
     begin
        $write("%c", `SOC_TOP.biu_pad_wdata[39:32]);
     end
     else if(cpu_wstrb[15:0] == 16'hf00)
     begin
        $write("%c", `SOC_TOP.biu_pad_wdata[71:64]);
     end
     else if(cpu_wstrb[15:0] == 16'hf000)
     begin
        $write("%c", `SOC_TOP.biu_pad_wdata[103:96]);
     end
    end
  end
  soc x_soc(
    .i_pad_clk           ( clk                  ),
    .i_pad_rst_b         ( rst_b                ),
    .biu_pad_htrans      (                      ),
    .biu_pad_hwrite      (                      ),
    .biu_pad_hwdata      (                      ),
    .biu_pad_haddr       (                      ),
    .prog_wen            ( 1'b0                 ),
    .prog_waddr          (                      ),
    .prog_wdata          (                      ),
    .uart2sys_en         ( 1'b0          ),
    .uart2sys_addr       ( uart2sys_addr[23:4]  ),
    .uart2sys_data       ( uart2sys_data        ),
    .sys_wren            ( 1'b0             ),
    .sys_data            ( sys_data             ),
    .sys_final_addr      ( sys_final_addr[23:4] ),
    .sysRAM_data         (                      ),
    .ram_wen             (                      )
  );
  int_mnt x_int_mnt(
  );
  
endmodule
